VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_32b_8192_1rw_freepdk45_sram_32x8192_1v
   CLASS BLOCK ;
   SIZE 444.4925 BY 762.6675 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  50.39 0.0 50.53 0.14 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  53.25 0.0 53.39 0.14 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  56.11 0.0 56.25 0.14 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  58.97 0.0 59.11 0.14 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  61.83 0.0 61.97 0.14 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  64.69 0.0 64.83 0.14 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  67.55 0.0 67.69 0.14 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  70.41 0.0 70.55 0.14 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  73.27 0.0 73.41 0.14 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  76.13 0.0 76.27 0.14 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  78.99 0.0 79.13 0.14 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  81.85 0.0 81.99 0.14 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  84.71 0.0 84.85 0.14 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  87.57 0.0 87.71 0.14 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  90.43 0.0 90.57 0.14 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  93.29 0.0 93.43 0.14 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  96.15 0.0 96.29 0.14 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  99.01 0.0 99.15 0.14 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  101.87 0.0 102.01 0.14 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  104.73 0.0 104.87 0.14 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  107.59 0.0 107.73 0.14 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  110.45 0.0 110.59 0.14 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  113.31 0.0 113.45 0.14 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  116.17 0.0 116.31 0.14 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  119.03 0.0 119.17 0.14 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  121.89 0.0 122.03 0.14 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  124.75 0.0 124.89 0.14 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  127.61 0.0 127.75 0.14 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  130.47 0.0 130.61 0.14 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  133.33 0.0 133.47 0.14 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  136.19 0.0 136.33 0.14 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  139.05 0.0 139.19 0.14 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  38.95 0.0 39.09 0.14 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  41.81 0.0 41.95 0.14 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  44.67 0.0 44.81 0.14 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER metal4 ;
         RECT  47.53 0.0 47.67 0.14 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 98.47 0.14 98.61 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 101.2 0.14 101.34 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 103.41 0.14 103.55 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 106.14 0.14 106.28 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 108.35 0.14 108.49 ;
      END
   END addr0[8]
   PIN addr0[9]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 111.08 0.14 111.22 ;
      END
   END addr0[9]
   PIN addr0[10]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 113.29 0.14 113.43 ;
      END
   END addr0[10]
   PIN addr0[11]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 116.02 0.14 116.16 ;
      END
   END addr0[11]
   PIN addr0[12]
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 118.23 0.14 118.37 ;
      END
   END addr0[12]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 37.37 0.14 37.51 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 40.1 0.14 40.24 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER metal3 ;
         RECT  0.0 37.605 0.14 37.745 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  78.2325 0.0 78.3725 0.14 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  89.62 0.0 89.76 0.14 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  101.1125 0.0 101.2525 0.14 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  112.415 0.0 112.555 0.14 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  123.695 0.0 123.835 0.14 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  134.975 0.0 135.115 0.14 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  146.255 0.0 146.395 0.14 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  157.535 0.0 157.675 0.14 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  168.815 0.0 168.955 0.14 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  180.095 0.0 180.235 0.14 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  191.375 0.0 191.515 0.14 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  202.655 0.0 202.795 0.14 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  213.935 0.0 214.075 0.14 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  225.215 0.0 225.355 0.14 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  236.495 0.0 236.635 0.14 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  247.775 0.0 247.915 0.14 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  259.055 0.0 259.195 0.14 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  270.335 0.0 270.475 0.14 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  281.615 0.0 281.755 0.14 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  292.895 0.0 293.035 0.14 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  304.175 0.0 304.315 0.14 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  315.455 0.0 315.595 0.14 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  326.735 0.0 326.875 0.14 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  338.015 0.0 338.155 0.14 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  349.295 0.0 349.435 0.14 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  360.575 0.0 360.715 0.14 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  371.855 0.0 371.995 0.14 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  383.135 0.0 383.275 0.14 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal4 ;
         RECT  394.415 0.0 394.555 0.14 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.3525 43.5025 444.4925 43.6425 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.3525 43.9725 444.4925 44.1125 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER metal3 ;
         RECT  444.3525 43.7375 444.4925 43.8775 ;
      END
   END dout0[31]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  0.0 0.0 0.7 762.6675 ;
         LAYER metal4 ;
         RECT  443.7925 0.0 444.4925 762.6675 ;
         LAYER metal3 ;
         RECT  0.0 761.9675 444.4925 762.6675 ;
         LAYER metal3 ;
         RECT  0.0 0.0 444.4925 0.7 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER metal4 ;
         RECT  442.3925 1.4 443.0925 761.2675 ;
         LAYER metal3 ;
         RECT  1.4 760.5675 443.0925 761.2675 ;
         LAYER metal4 ;
         RECT  1.4 1.4 2.1 761.2675 ;
         LAYER metal3 ;
         RECT  1.4 1.4 443.0925 2.1 ;
      END
   END gnd
   OBS
   LAYER  metal1 ;
      RECT  0.14 0.14 444.3525 762.5275 ;
   LAYER  metal2 ;
      RECT  0.14 0.14 444.3525 762.5275 ;
   LAYER  metal3 ;
      RECT  0.28 98.33 444.3525 98.75 ;
      RECT  0.14 98.75 0.28 101.06 ;
      RECT  0.14 101.48 0.28 103.27 ;
      RECT  0.14 103.69 0.28 106.0 ;
      RECT  0.14 106.42 0.28 108.21 ;
      RECT  0.14 108.63 0.28 110.94 ;
      RECT  0.14 111.36 0.28 113.15 ;
      RECT  0.14 113.57 0.28 115.88 ;
      RECT  0.14 116.3 0.28 118.09 ;
      RECT  0.14 40.38 0.28 98.33 ;
      RECT  0.14 37.885 0.28 39.96 ;
      RECT  0.28 43.3625 444.2125 43.7825 ;
      RECT  0.28 43.7825 444.2125 98.33 ;
      RECT  444.2125 44.2525 444.3525 98.33 ;
      RECT  0.14 118.51 0.28 761.8275 ;
      RECT  0.14 0.84 0.28 37.23 ;
      RECT  444.2125 0.84 444.3525 43.3625 ;
      RECT  0.28 98.75 1.26 760.4275 ;
      RECT  0.28 760.4275 1.26 761.4075 ;
      RECT  0.28 761.4075 1.26 761.8275 ;
      RECT  1.26 98.75 443.2325 760.4275 ;
      RECT  1.26 761.4075 443.2325 761.8275 ;
      RECT  443.2325 98.75 444.3525 760.4275 ;
      RECT  443.2325 760.4275 444.3525 761.4075 ;
      RECT  443.2325 761.4075 444.3525 761.8275 ;
      RECT  0.28 0.84 1.26 1.26 ;
      RECT  0.28 1.26 1.26 2.24 ;
      RECT  0.28 2.24 1.26 43.3625 ;
      RECT  1.26 0.84 443.2325 1.26 ;
      RECT  1.26 2.24 443.2325 43.3625 ;
      RECT  443.2325 0.84 444.2125 1.26 ;
      RECT  443.2325 1.26 444.2125 2.24 ;
      RECT  443.2325 2.24 444.2125 43.3625 ;
   LAYER  metal4 ;
      RECT  50.11 0.42 50.81 762.5275 ;
      RECT  50.81 0.14 52.97 0.42 ;
      RECT  53.67 0.14 55.83 0.42 ;
      RECT  56.53 0.14 58.69 0.42 ;
      RECT  59.39 0.14 61.55 0.42 ;
      RECT  62.25 0.14 64.41 0.42 ;
      RECT  65.11 0.14 67.27 0.42 ;
      RECT  67.97 0.14 70.13 0.42 ;
      RECT  70.83 0.14 72.99 0.42 ;
      RECT  73.69 0.14 75.85 0.42 ;
      RECT  79.41 0.14 81.57 0.42 ;
      RECT  82.27 0.14 84.43 0.42 ;
      RECT  85.13 0.14 87.29 0.42 ;
      RECT  90.85 0.14 93.01 0.42 ;
      RECT  93.71 0.14 95.87 0.42 ;
      RECT  96.57 0.14 98.73 0.42 ;
      RECT  102.29 0.14 104.45 0.42 ;
      RECT  105.15 0.14 107.31 0.42 ;
      RECT  108.01 0.14 110.17 0.42 ;
      RECT  113.73 0.14 115.89 0.42 ;
      RECT  116.59 0.14 118.75 0.42 ;
      RECT  119.45 0.14 121.61 0.42 ;
      RECT  125.17 0.14 127.33 0.42 ;
      RECT  128.03 0.14 130.19 0.42 ;
      RECT  130.89 0.14 133.05 0.42 ;
      RECT  136.61 0.14 138.77 0.42 ;
      RECT  39.37 0.14 41.53 0.42 ;
      RECT  42.23 0.14 44.39 0.42 ;
      RECT  45.09 0.14 47.25 0.42 ;
      RECT  47.95 0.14 50.11 0.42 ;
      RECT  76.55 0.14 77.9525 0.42 ;
      RECT  78.6525 0.14 78.71 0.42 ;
      RECT  87.99 0.14 89.34 0.42 ;
      RECT  90.04 0.14 90.15 0.42 ;
      RECT  99.43 0.14 100.8325 0.42 ;
      RECT  101.5325 0.14 101.59 0.42 ;
      RECT  110.87 0.14 112.135 0.42 ;
      RECT  112.835 0.14 113.03 0.42 ;
      RECT  122.31 0.14 123.415 0.42 ;
      RECT  124.115 0.14 124.47 0.42 ;
      RECT  133.75 0.14 134.695 0.42 ;
      RECT  135.395 0.14 135.91 0.42 ;
      RECT  139.47 0.14 145.975 0.42 ;
      RECT  146.675 0.14 157.255 0.42 ;
      RECT  157.955 0.14 168.535 0.42 ;
      RECT  169.235 0.14 179.815 0.42 ;
      RECT  180.515 0.14 191.095 0.42 ;
      RECT  191.795 0.14 202.375 0.42 ;
      RECT  203.075 0.14 213.655 0.42 ;
      RECT  214.355 0.14 224.935 0.42 ;
      RECT  225.635 0.14 236.215 0.42 ;
      RECT  236.915 0.14 247.495 0.42 ;
      RECT  248.195 0.14 258.775 0.42 ;
      RECT  259.475 0.14 270.055 0.42 ;
      RECT  270.755 0.14 281.335 0.42 ;
      RECT  282.035 0.14 292.615 0.42 ;
      RECT  293.315 0.14 303.895 0.42 ;
      RECT  304.595 0.14 315.175 0.42 ;
      RECT  315.875 0.14 326.455 0.42 ;
      RECT  327.155 0.14 337.735 0.42 ;
      RECT  338.435 0.14 349.015 0.42 ;
      RECT  349.715 0.14 360.295 0.42 ;
      RECT  360.995 0.14 371.575 0.42 ;
      RECT  372.275 0.14 382.855 0.42 ;
      RECT  383.555 0.14 394.135 0.42 ;
      RECT  0.98 0.14 38.67 0.42 ;
      RECT  394.835 0.14 443.5125 0.42 ;
      RECT  50.81 0.42 442.1125 1.12 ;
      RECT  50.81 1.12 442.1125 761.5475 ;
      RECT  50.81 761.5475 442.1125 762.5275 ;
      RECT  442.1125 0.42 443.3725 1.12 ;
      RECT  442.1125 761.5475 443.3725 762.5275 ;
      RECT  443.3725 0.42 443.5125 1.12 ;
      RECT  443.3725 1.12 443.5125 761.5475 ;
      RECT  443.3725 761.5475 443.5125 762.5275 ;
      RECT  0.98 0.42 1.12 1.12 ;
      RECT  0.98 1.12 1.12 761.5475 ;
      RECT  0.98 761.5475 1.12 762.5275 ;
      RECT  1.12 0.42 2.38 1.12 ;
      RECT  1.12 761.5475 2.38 762.5275 ;
      RECT  2.38 0.42 50.11 1.12 ;
      RECT  2.38 1.12 50.11 761.5475 ;
      RECT  2.38 761.5475 50.11 762.5275 ;
   END
END    sram_32b_8192_1rw_freepdk45_sram_32x8192_1v
END    LIBRARY
